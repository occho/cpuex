library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;

entity prom is

	port (
		clka : in std_logic;
		addra : in std_logic_vector(11 downto 0);
		douta : out std_logic_vector(31 downto 0));

end prom;

architecture RTL of prom is
	subtype word_t is std_logic_vector(31 downto 0);
	type mem_t is array (0 to 4095) of word_t;
	signal addr_in	: integer range 0 to 4095;

	constant mem : mem_t := (
x"0000004c",
x"00000000",
x"3f800000",
x"bf800000",
x"00800000",
x"4b000000",
x"4b000000",
x"41400000",
x"41300000",
x"41200000",
x"41100000",
x"41000000",
x"40e00000",
x"40c00000",
x"40a00000",
x"40800000",
x"40400000",
x"3f800000",
x"00000000",
x"40000000",
x"a0000000",
x"080001d3",
x"a0000000",
x"a0000000",
x"a0630002",
x"a0000000",
x"a0000000",
x"00622820",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"68a2000e",
x"a0000000",
x"a0000000",
x"28a2000b",
x"a0000000",
x"a0000000",
x"ac440000",
x"a0000000",
x"a0000000",
x"20420004",
x"a0000000",
x"a0000000",
x"08000020",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0630002",
x"a0000000",
x"a0000000",
x"00622020",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"6882000e",
x"a0000000",
x"a0000000",
x"2882000b",
x"a0000000",
x"a0000000",
x"e4400000",
x"a0000000",
x"a0000000",
x"20420004",
x"a0000000",
x"a0000000",
x"0800003b",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"c4640000",
x"a0000000",
x"a0000000",
x"e880003e",
x"a0000000",
x"a0000000",
x"c880003b",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"20030010",
x"a0000000",
x"a0000000",
x"c4620000",
x"a0000000",
x"a0000000",
x"e802000b",
x"a0000000",
x"a0000000",
x"c8020008",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"44200807",
x"a0000000",
x"a0000000",
x"e8200050",
x"a0000000",
x"a0000000",
x"c820004d",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"20030004",
x"a0000000",
x"a0000000",
x"c4630000",
x"a0000000",
x"a0000000",
x"44030000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20030010",
x"a0000000",
x"a0000000",
x"c4620000",
x"a0000000",
x"a0000000",
x"e8020008",
x"a0000000",
x"a0000000",
x"c8020005",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"e801000e",
x"a0000000",
x"a0000000",
x"c801000b",
x"a0000000",
x"a0000000",
x"20030004",
x"a0000000",
x"a0000000",
x"c4630000",
x"a0000000",
x"a0000000",
x"44030001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"c000004d",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"68030011",
x"a0000000",
x"a0000000",
x"2803000e",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"c00000ef",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20050010",
x"a0000000",
x"a0000000",
x"c4a10000",
x"a0000000",
x"a0000000",
x"20050014",
x"a0000000",
x"a0000000",
x"8ca40000",
x"a0000000",
x"a0000000",
x"2005000c",
x"a0000000",
x"a0000000",
x"8ca50000",
x"a0000000",
x"a0000000",
x"68a30014",
x"a0000000",
x"a0000000",
x"28a30011",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"44010001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"c4820000",
x"a0000000",
x"a0000000",
x"00651822",
x"a0000000",
x"a0000000",
x"44411000",
x"a0000000",
x"a0000000",
x"68a3fff9",
x"a0000000",
x"a0000000",
x"28a3fff6",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"44010001",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"c4610000",
x"a0000000",
x"a0000000",
x"e8200011",
x"a0000000",
x"a0000000",
x"c820000e",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"c0000152",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"c000004d",
x"a0000000",
x"a0000000",
x"20040010",
x"a0000000",
x"a0000000",
x"c4820000",
x"a0000000",
x"a0000000",
x"20040014",
x"a0000000",
x"a0000000",
x"8c840000",
x"a0000000",
x"a0000000",
x"e8400014",
x"a0000000",
x"a0000000",
x"c8400011",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c230000",
x"a0000000",
x"a0000000",
x"00641822",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"2005000c",
x"a0000000",
x"a0000000",
x"8ca50000",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"00651820",
x"a0000000",
x"a0000000",
x"e840fff9",
x"a0000000",
x"a0000000",
x"c840fff6",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c250000",
x"a0000000",
x"a0000000",
x"00a42822",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"0800013a",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"c00001a0",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"203f0000",
x"a0000000",
x"a0000000",
x"40210030",
x"a0000000",
x"a0000000",
x"201c0001",
x"a0000000",
x"a0000000",
x"201dffff",
x"a0000000",
x"a0000000",
x"201b0044",
x"a0000000",
x"a0000000",
x"c7700000",
x"a0000000",
x"a0000000",
x"201b0024",
x"a0000000",
x"a0000000",
x"c7710000",
x"a0000000",
x"a0000000",
x"201b0028",
x"a0000000",
x"a0000000",
x"c7720000",
x"a0000000",
x"a0000000",
x"201b002c",
x"a0000000",
x"a0000000",
x"c7730000",
x"a0000000",
x"a0000000",
x"201b0030",
x"a0000000",
x"a0000000",
x"c7740000",
x"a0000000",
x"a0000000",
x"201b0034",
x"a0000000",
x"a0000000",
x"c7750000",
x"a0000000",
x"a0000000",
x"201b0038",
x"a0000000",
x"a0000000",
x"c7760000",
x"a0000000",
x"a0000000",
x"201b003c",
x"a0000000",
x"a0000000",
x"c7770000",
x"a0000000",
x"a0000000",
x"201b0040",
x"a0000000",
x"a0000000",
x"c7780000",
x"a0000000",
x"a0000000",
x"201b0048",
x"a0000000",
x"a0000000",
x"c7790000",
x"a0000000",
x"a0000000",
x"201b0018",
x"a0000000",
x"a0000000",
x"c77a0000",
x"a0000000",
x"a0000000",
x"201b001c",
x"a0000000",
x"a0000000",
x"c77b0000",
x"a0000000",
x"a0000000",
x"201b0020",
x"a0000000",
x"a0000000",
x"c77c0000",
x"a0000000",
x"a0000000",
x"47200006",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e20004",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e20008",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e2000c",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e20010",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040001",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e20014",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e20018",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"46000006",
x"a0000000",
x"a0000000",
x"afe2002c",
x"a0000000",
x"a0000000",
x"43e2001c",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000032",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"8fe2002c",
x"a0000000",
x"a0000000",
x"20030002",
x"a0000000",
x"a0000000",
x"20040003",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000895",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"afe30020",
x"a0000000",
x"a0000000",
x"20040003",
x"a0000000",
x"a0000000",
x"20050002",
x"a0000000",
x"a0000000",
x"ac230004",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"20a40000",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"c0000895",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"afe30024",
x"a0000000",
x"a0000000",
x"20040002",
x"a0000000",
x"a0000000",
x"20050002",
x"a0000000",
x"a0000000",
x"ac230008",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"20a40000",
x"a0000000",
x"a0000000",
x"40210010",
x"a0000000",
x"a0000000",
x"c0000895",
x"a0000000",
x"a0000000",
x"20210010",
x"a0000000",
x"a0000000",
x"20680000",
x"a0000000",
x"a0000000",
x"afe80028",
x"a0000000",
x"a0000000",
x"8c260004",
x"a0000000",
x"a0000000",
x"8cc30000",
x"a0000000",
x"a0000000",
x"47000006",
x"a0000000",
x"a0000000",
x"e4600000",
x"a0000000",
x"a0000000",
x"8cc30000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"e460fffc",
x"a0000000",
x"a0000000",
x"8cc30000",
x"a0000000",
x"a0000000",
x"46e00006",
x"a0000000",
x"a0000000",
x"e460fff8",
x"a0000000",
x"a0000000",
x"8cc3fffc",
x"a0000000",
x"a0000000",
x"46c00006",
x"a0000000",
x"a0000000",
x"e4600000",
x"a0000000",
x"a0000000",
x"8cc3fffc",
x"a0000000",
x"a0000000",
x"46a00006",
x"a0000000",
x"a0000000",
x"e460fffc",
x"a0000000",
x"a0000000",
x"8cc3fffc",
x"a0000000",
x"a0000000",
x"46800006",
x"a0000000",
x"a0000000",
x"e460fff8",
x"a0000000",
x"a0000000",
x"8c270008",
x"a0000000",
x"a0000000",
x"8ce30000",
x"a0000000",
x"a0000000",
x"46600006",
x"a0000000",
x"a0000000",
x"e4600000",
x"a0000000",
x"a0000000",
x"8ce30000",
x"a0000000",
x"a0000000",
x"46400006",
x"a0000000",
x"a0000000",
x"e460fffc",
x"a0000000",
x"a0000000",
x"8ce3fffc",
x"a0000000",
x"a0000000",
x"46200006",
x"a0000000",
x"a0000000",
x"e4600000",
x"a0000000",
x"a0000000",
x"8ce3fffc",
x"a0000000",
x"a0000000",
x"47800006",
x"a0000000",
x"a0000000",
x"e460fffc",
x"a0000000",
x"a0000000",
x"8ce3fff8",
x"a0000000",
x"a0000000",
x"47600006",
x"a0000000",
x"a0000000",
x"e4600000",
x"a0000000",
x"a0000000",
x"8ce3fff8",
x"a0000000",
x"a0000000",
x"47400006",
x"a0000000",
x"a0000000",
x"e460fffc",
x"a0000000",
x"a0000000",
x"20030002",
x"a0000000",
x"a0000000",
x"20040003",
x"a0000000",
x"a0000000",
x"20050002",
x"a0000000",
x"a0000000",
x"ac28000c",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c0000835",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"8c23000c",
x"a0000000",
x"a0000000",
x"8c640000",
x"a0000000",
x"a0000000",
x"c4800000",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000019d",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000047b",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"ac230014",
x"a0000000",
x"a0000000",
x"2003000a",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"8c230014",
x"a0000000",
x"a0000000",
x"8c23000c",
x"a0000000",
x"a0000000",
x"8c640000",
x"a0000000",
x"a0000000",
x"c480fffc",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000019d",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000047b",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"ac230014",
x"a0000000",
x"a0000000",
x"2003000a",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"8c230014",
x"a0000000",
x"a0000000",
x"8c23000c",
x"a0000000",
x"a0000000",
x"8c64fffc",
x"a0000000",
x"a0000000",
x"c4800000",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000019d",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000047b",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"ac230014",
x"a0000000",
x"a0000000",
x"2003000a",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"8c230014",
x"a0000000",
x"a0000000",
x"8c23000c",
x"a0000000",
x"a0000000",
x"8c63fffc",
x"a0000000",
x"a0000000",
x"c460fffc",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000019d",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c000047b",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"ac230014",
x"a0000000",
x"a0000000",
x"2003000a",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"8c230014",
x"a0000000",
x"a0000000",
x"0800044a",
x"0800044a",
x"0800044a",
x"a0000000",
x"a0000000",
x"00a63820",
x"a0000000",
x"a0000000",
x"a8e70001",
x"a0000000",
x"a0000000",
x"00e44018",
x"a0000000",
x"a0000000",
x"00c54822",
x"a0000000",
x"a0000000",
x"6b890008",
x"a0000000",
x"a0000000",
x"20a30000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"69030011",
x"a0000000",
x"a0000000",
x"49030008",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20e60000",
x"a0000000",
x"a0000000",
x"0800044e",
x"a0000000",
x"a0000000",
x"20e50000",
x"a0000000",
x"a0000000",
x"0800044e",
x"a0000000",
x"a0000000",
x"686002a5",
x"a0000000",
x"a0000000",
x"3c8005f5",
x"a0000000",
x"a0000000",
x"1c80e100",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"20060003",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"3c8005f5",
x"a0000000",
x"a0000000",
x"1c80e100",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c250000",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac240004",
x"a0000000",
x"a0000000",
x"68030008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"080004bd",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"3c800098",
x"a0000000",
x"a0000000",
x"1c809680",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c270004",
x"a0000000",
x"a0000000",
x"ac230008",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210010",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210010",
x"a0000000",
x"a0000000",
x"3c800098",
x"a0000000",
x"a0000000",
x"1c809680",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c250004",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac24000c",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250008",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"08000508",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"08000517",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"3c80000f",
x"a0000000",
x"a0000000",
x"1c804240",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c27000c",
x"a0000000",
x"a0000000",
x"ac230010",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210018",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210018",
x"a0000000",
x"a0000000",
x"3c80000f",
x"a0000000",
x"a0000000",
x"1c804240",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c25000c",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac240014",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250010",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"08000562",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"08000571",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"3c800001",
x"a0000000",
x"a0000000",
x"1c8086a0",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c270014",
x"a0000000",
x"a0000000",
x"ac230018",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210020",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210020",
x"a0000000",
x"a0000000",
x"3c800001",
x"a0000000",
x"a0000000",
x"1c8086a0",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c250014",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac24001c",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250018",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"080005bc",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"080005cb",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20042710",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c27001c",
x"a0000000",
x"a0000000",
x"ac230020",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210028",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210028",
x"a0000000",
x"a0000000",
x"20042710",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c25001c",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac240024",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250020",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"08000610",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"0800061f",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"200403e8",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c270024",
x"a0000000",
x"a0000000",
x"ac230028",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210030",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210030",
x"a0000000",
x"a0000000",
x"606403e8",
x"a0000000",
x"a0000000",
x"8c250024",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac24002c",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250028",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"08000661",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"08000670",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040064",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c27002c",
x"a0000000",
x"a0000000",
x"ac230030",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210038",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210038",
x"a0000000",
x"a0000000",
x"60640064",
x"a0000000",
x"a0000000",
x"8c25002c",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac240034",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250030",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"080006b2",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"080006c1",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"2004000a",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"8c270034",
x"a0000000",
x"a0000000",
x"ac230038",
x"a0000000",
x"a0000000",
x"20e30000",
x"a0000000",
x"a0000000",
x"40210040",
x"a0000000",
x"a0000000",
x"c000044e",
x"a0000000",
x"a0000000",
x"20210040",
x"a0000000",
x"a0000000",
x"6064000a",
x"a0000000",
x"a0000000",
x"8c250034",
x"a0000000",
x"a0000000",
x"00a42022",
x"a0000000",
x"a0000000",
x"ac24003c",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"8c250038",
x"a0000000",
x"a0000000",
x"48a00008",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"08000703",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"08000712",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20030030",
x"a0000000",
x"a0000000",
x"8c24003c",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"2004002d",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"04800001",
x"a0000000",
x"a0000000",
x"8c230000",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"0800047b",
x"a0000000",
x"a0000000",
x"8fc4ffec",
x"a0000000",
x"a0000000",
x"8fc5fff0",
x"a0000000",
x"a0000000",
x"8fc6fff4",
x"a0000000",
x"a0000000",
x"8fc7fff8",
x"a0000000",
x"a0000000",
x"8fc8fffc",
x"a0000000",
x"a0000000",
x"6860003b",
x"a0000000",
x"a0000000",
x"a0a90002",
x"a0000000",
x"a0000000",
x"4cc93000",
x"a0000000",
x"a0000000",
x"a0890002",
x"a0000000",
x"a0000000",
x"00c90031",
x"a0000000",
x"a0000000",
x"a0a50002",
x"a0000000",
x"a0000000",
x"4d052800",
x"a0000000",
x"a0000000",
x"a0680002",
x"a0000000",
x"a0000000",
x"00a80831",
x"a0000000",
x"a0000000",
x"a0650002",
x"a0000000",
x"a0000000",
x"4ce52800",
x"a0000000",
x"a0000000",
x"a0870002",
x"a0000000",
x"a0000000",
x"00a71031",
x"a0000000",
x"a0000000",
x"44220802",
x"a0000000",
x"a0000000",
x"44010000",
x"a0000000",
x"a0000000",
x"a0840002",
x"a0000000",
x"a0000000",
x"00c40039",
x"a0000000",
x"a0000000",
x"40630001",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"03600008",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"8fc4ffec",
x"a0000000",
x"a0000000",
x"8fc5fff0",
x"a0000000",
x"a0000000",
x"8fc6fff4",
x"a0000000",
x"a0000000",
x"8fc7fff8",
x"a0000000",
x"a0000000",
x"8fc8fffc",
x"a0000000",
x"a0000000",
x"68600047",
x"a0000000",
x"a0000000",
x"20490000",
x"a0000000",
x"a0000000",
x"20420018",
x"a0000000",
x"a0000000",
x"200a0733",
x"a0000000",
x"a0000000",
x"ad2a0000",
x"a0000000",
x"a0000000",
x"ad23ffec",
x"a0000000",
x"a0000000",
x"ad25fff0",
x"a0000000",
x"a0000000",
x"ad26fff4",
x"a0000000",
x"a0000000",
x"ad27fff8",
x"a0000000",
x"a0000000",
x"ad28fffc",
x"a0000000",
x"a0000000",
x"40840001",
x"a0000000",
x"a0000000",
x"ac3e0000",
x"a0000000",
x"a0000000",
x"ac230004",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"213e0000",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"03600030",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"8c230004",
x"a0000000",
x"a0000000",
x"40630001",
x"a0000000",
x"a0000000",
x"8c3e0000",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"03600008",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"8fc4ffec",
x"a0000000",
x"a0000000",
x"8fc5fff0",
x"a0000000",
x"a0000000",
x"8fc6fff4",
x"a0000000",
x"a0000000",
x"8fc7fff8",
x"a0000000",
x"a0000000",
x"8fc8fffc",
x"a0000000",
x"a0000000",
x"68600047",
x"a0000000",
x"a0000000",
x"20490000",
x"a0000000",
x"a0000000",
x"20420018",
x"a0000000",
x"a0000000",
x"200a0781",
x"a0000000",
x"a0000000",
x"ad2a0000",
x"a0000000",
x"a0000000",
x"ad25ffec",
x"a0000000",
x"a0000000",
x"ad23fff0",
x"a0000000",
x"a0000000",
x"ad26fff4",
x"a0000000",
x"a0000000",
x"ad27fff8",
x"a0000000",
x"a0000000",
x"ad28fffc",
x"a0000000",
x"a0000000",
x"40840001",
x"a0000000",
x"a0000000",
x"ac3e0000",
x"a0000000",
x"a0000000",
x"ac230004",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"213e0000",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"03600030",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"8c230004",
x"a0000000",
x"a0000000",
x"40630001",
x"a0000000",
x"a0000000",
x"8c3e0000",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"03600008",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"205e0000",
x"a0000000",
x"a0000000",
x"20420018",
x"a0000000",
x"a0000000",
x"200907db",
x"a0000000",
x"a0000000",
x"afc90000",
x"a0000000",
x"a0000000",
x"afc5ffec",
x"a0000000",
x"a0000000",
x"afc4fff0",
x"a0000000",
x"a0000000",
x"afc8fff4",
x"a0000000",
x"a0000000",
x"afc7fff8",
x"a0000000",
x"a0000000",
x"afc6fffc",
x"a0000000",
x"a0000000",
x"40630001",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"03600008",
x"a0000000",
x"a0000000",
x"8fc4fff8",
x"a0000000",
x"a0000000",
x"8fc5fffc",
x"a0000000",
x"a0000000",
x"68600032",
x"a0000000",
x"a0000000",
x"46000006",
x"a0000000",
x"a0000000",
x"ac3e0000",
x"a0000000",
x"a0000000",
x"ac250004",
x"a0000000",
x"a0000000",
x"ac230008",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"40210010",
x"a0000000",
x"a0000000",
x"c0000032",
x"a0000000",
x"a0000000",
x"20210010",
x"a0000000",
x"a0000000",
x"8c240008",
x"a0000000",
x"a0000000",
x"a0850002",
x"a0000000",
x"a0000000",
x"8c260004",
x"a0000000",
x"a0000000",
x"6cc51800",
x"a0000000",
x"a0000000",
x"40830001",
x"a0000000",
x"a0000000",
x"8c3e0000",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"03600008",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"43e5001c",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"ac240004",
x"a0000000",
x"a0000000",
x"20a40000",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"c0000017",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"205e0000",
x"a0000000",
x"a0000000",
x"2042000c",
x"a0000000",
x"a0000000",
x"20040859",
x"a0000000",
x"a0000000",
x"afc40000",
x"a0000000",
x"a0000000",
x"8c240004",
x"a0000000",
x"a0000000",
x"afc4fff8",
x"a0000000",
x"a0000000",
x"afc3fffc",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"40840001",
x"a0000000",
x"a0000000",
x"ac230008",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"8fdb0000",
x"a0000000",
x"a0000000",
x"40210010",
x"a0000000",
x"a0000000",
x"03600030",
x"a0000000",
x"a0000000",
x"20210010",
x"a0000000",
x"a0000000",
x"8c230008",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000"
	 );


begin
	prom_sim: process(clka)
	begin
		if rising_edge(clka) then
			addr_in <= conv_integer(addra);
			douta <= mem(addr_in);
		end if;
	end process;

end RTL;



