library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;

entity prom is

	port (
		clka : in std_logic;
		addra : in std_logic_vector(11 downto 0);
		douta : out std_logic_vector(31 downto 0));

end prom;

architecture RTL of prom is
	subtype word_t is std_logic_vector(31 downto 0);
	type mem_t is array (0 to 4095) of word_t;
	signal addr_in	: integer range 0 to 4095;

	constant mem : mem_t := (
x"00000034",
x"00000000",
x"3f800000",
x"bf800000",
x"00800000",
x"4b000000",
x"4b000000",
x"40c00000",
x"40a00000",
x"40800000",
x"40400000",
x"3f800000",
x"49742400",
x"40000000",
x"a0000000",
x"080001cd",
x"a0000000",
x"a0000000",
x"a0630002",
x"a0000000",
x"a0000000",
x"00622820",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"68a2000e",
x"a0000000",
x"a0000000",
x"28a2000b",
x"a0000000",
x"a0000000",
x"ac440000",
x"a0000000",
x"a0000000",
x"20420004",
x"a0000000",
x"a0000000",
x"0800001a",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0630002",
x"a0000000",
x"a0000000",
x"00622020",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"6882000e",
x"a0000000",
x"a0000000",
x"2882000b",
x"a0000000",
x"a0000000",
x"e4400000",
x"a0000000",
x"a0000000",
x"20420004",
x"a0000000",
x"a0000000",
x"08000035",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"c4640000",
x"a0000000",
x"a0000000",
x"e880003e",
x"a0000000",
x"a0000000",
x"c880003b",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"20030010",
x"a0000000",
x"a0000000",
x"c4620000",
x"a0000000",
x"a0000000",
x"e802000b",
x"a0000000",
x"a0000000",
x"c8020008",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"44200807",
x"a0000000",
x"a0000000",
x"e8200050",
x"a0000000",
x"a0000000",
x"c820004d",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"20030004",
x"a0000000",
x"a0000000",
x"c4630000",
x"a0000000",
x"a0000000",
x"44030000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20030010",
x"a0000000",
x"a0000000",
x"c4620000",
x"a0000000",
x"a0000000",
x"e8020008",
x"a0000000",
x"a0000000",
x"c8020005",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"e801000e",
x"a0000000",
x"a0000000",
x"c801000b",
x"a0000000",
x"a0000000",
x"20030004",
x"a0000000",
x"a0000000",
x"c4630000",
x"a0000000",
x"a0000000",
x"44030001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"c0000047",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"68030011",
x"a0000000",
x"a0000000",
x"2803000e",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"c00000e9",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20050010",
x"a0000000",
x"a0000000",
x"c4a10000",
x"a0000000",
x"a0000000",
x"20050014",
x"a0000000",
x"a0000000",
x"8ca40000",
x"a0000000",
x"a0000000",
x"2005000c",
x"a0000000",
x"a0000000",
x"8ca50000",
x"a0000000",
x"a0000000",
x"68a30014",
x"a0000000",
x"a0000000",
x"28a30011",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"44010001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"c4820000",
x"a0000000",
x"a0000000",
x"00651822",
x"a0000000",
x"a0000000",
x"44411000",
x"a0000000",
x"a0000000",
x"68a3fff9",
x"a0000000",
x"a0000000",
x"28a3fff6",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"44010001",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"c4610000",
x"a0000000",
x"a0000000",
x"e8200011",
x"a0000000",
x"a0000000",
x"c820000e",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"c000014c",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"c0000047",
x"a0000000",
x"a0000000",
x"20040010",
x"a0000000",
x"a0000000",
x"c4820000",
x"a0000000",
x"a0000000",
x"20040014",
x"a0000000",
x"a0000000",
x"8c840000",
x"a0000000",
x"a0000000",
x"e8400014",
x"a0000000",
x"a0000000",
x"c8400011",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c230000",
x"a0000000",
x"a0000000",
x"00641822",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"2005000c",
x"a0000000",
x"a0000000",
x"8ca50000",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"00651820",
x"a0000000",
x"a0000000",
x"e840fff9",
x"a0000000",
x"a0000000",
x"c840fff6",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c250000",
x"a0000000",
x"a0000000",
x"00a42822",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"08000134",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"c000019a",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"203f0000",
x"a0000000",
x"a0000000",
x"40210020",
x"a0000000",
x"a0000000",
x"201c0001",
x"a0000000",
x"a0000000",
x"201dffff",
x"a0000000",
x"a0000000",
x"201b0018",
x"a0000000",
x"a0000000",
x"c7700000",
x"a0000000",
x"a0000000",
x"201b001c",
x"a0000000",
x"a0000000",
x"c7710000",
x"a0000000",
x"a0000000",
x"201b0020",
x"a0000000",
x"a0000000",
x"c7720000",
x"a0000000",
x"a0000000",
x"201b0024",
x"a0000000",
x"a0000000",
x"c7730000",
x"a0000000",
x"a0000000",
x"201b0028",
x"a0000000",
x"a0000000",
x"c7740000",
x"a0000000",
x"a0000000",
x"201b002c",
x"a0000000",
x"a0000000",
x"c7750000",
x"a0000000",
x"a0000000",
x"201b0030",
x"a0000000",
x"a0000000",
x"c7760000",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20004",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000011",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20008",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000011",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e2000c",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000011",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20010",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000011",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040001",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20014",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000011",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20018",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000011",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20440000",
x"a0000000",
x"a0000000",
x"2042000c",
x"a0000000",
x"a0000000",
x"e493fff8",
x"a0000000",
x"a0000000",
x"e496fffc",
x"a0000000",
x"a0000000",
x"e4940000",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"2042000c",
x"a0000000",
x"a0000000",
x"e470fff8",
x"a0000000",
x"a0000000",
x"e471fffc",
x"a0000000",
x"a0000000",
x"e4720000",
x"a0000000",
x"a0000000",
x"20850000",
x"a0000000",
x"a0000000",
x"20640000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000574",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"46a00002",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000197",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"20680000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c000030a",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"080002d9",
x"080002d9",
x"080002d9",
x"a0000000",
x"a0000000",
x"00a61820",
x"a0000000",
x"a0000000",
x"a8640001",
x"a0000000",
x"a0000000",
x"00874818",
x"a0000000",
x"a0000000",
x"00c51822",
x"a0000000",
x"a0000000",
x"6b830008",
x"a0000000",
x"a0000000",
x"20a30000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"69280011",
x"a0000000",
x"a0000000",
x"49280008",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20860000",
x"a0000000",
x"a0000000",
x"080002dd",
x"a0000000",
x"a0000000",
x"20850000",
x"a0000000",
x"a0000000",
x"080002dd",
x"a0000000",
x"a0000000",
x"6900024b",
x"a0000000",
x"a0000000",
x"3ce005f5",
x"a0000000",
x"a0000000",
x"1ce0e100",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"20060003",
x"a0000000",
x"a0000000",
x"ac280000",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"3c8005f5",
x"a0000000",
x"a0000000",
x"1c80e100",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280000",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"68030008",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"08000349",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"3ce00098",
x"a0000000",
x"a0000000",
x"1ce09680",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280004",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"3c800098",
x"a0000000",
x"a0000000",
x"1c809680",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280004",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49400008",
x"a0000000",
x"a0000000",
x"200b0000",
x"a0000000",
x"a0000000",
x"08000388",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"08000397",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"3ce0000f",
x"a0000000",
x"a0000000",
x"1ce04240",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280008",
x"a0000000",
x"a0000000",
x"40210010",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"20210010",
x"a0000000",
x"a0000000",
x"3c80000f",
x"a0000000",
x"a0000000",
x"1c804240",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280008",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49600008",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"080003d6",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"080003e5",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"3ce00001",
x"a0000000",
x"a0000000",
x"1ce086a0",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac28000c",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"3c800001",
x"a0000000",
x"a0000000",
x"1c8086a0",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c28000c",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49400008",
x"a0000000",
x"a0000000",
x"200b0000",
x"a0000000",
x"a0000000",
x"08000424",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"08000433",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"20072710",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280010",
x"a0000000",
x"a0000000",
x"40210018",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"20210018",
x"a0000000",
x"a0000000",
x"20042710",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280010",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49600008",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"0800046c",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"0800047b",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"200703e8",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280014",
x"a0000000",
x"a0000000",
x"4021001c",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"2021001c",
x"a0000000",
x"a0000000",
x"606403e8",
x"a0000000",
x"a0000000",
x"8c280014",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49400008",
x"a0000000",
x"a0000000",
x"200b0000",
x"a0000000",
x"a0000000",
x"080004b1",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"080004c0",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"20070064",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280018",
x"a0000000",
x"a0000000",
x"40210020",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"20210020",
x"a0000000",
x"a0000000",
x"60640064",
x"a0000000",
x"a0000000",
x"8c280018",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49600008",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"080004f6",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"08000505",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"2007000a",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac28001c",
x"a0000000",
x"a0000000",
x"40210024",
x"a0000000",
x"a0000000",
x"c00002dd",
x"a0000000",
x"a0000000",
x"20210024",
x"a0000000",
x"a0000000",
x"6064000a",
x"a0000000",
x"a0000000",
x"8c28001c",
x"a0000000",
x"a0000000",
x"01042022",
x"a0000000",
x"a0000000",
x"6803001a",
x"a0000000",
x"a0000000",
x"49400008",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"0800053b",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20050001",
x"a0000000",
x"a0000000",
x"0800054a",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20050001",
x"a0000000",
x"a0000000",
x"20030030",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"2003002d",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"00084022",
x"a0000000",
x"a0000000",
x"0800030a",
x"a0000000",
x"a0000000",
x"c4600000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"c460fffc",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"c460fff8",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"20a30000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000562",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000562",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"44201002",
x"a0000000",
x"a0000000",
x"20a30000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000568",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c0000568",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"44200002",
x"a0000000",
x"a0000000",
x"44401000",
x"a0000000",
x"a0000000",
x"20a30000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c000056e",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c000056e",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"44200002",
x"a0000000",
x"a0000000",
x"44400000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000"
	 );


begin
	prom_sim: process(clka)
	begin
		if rising_edge(clka) then
			addr_in <= conv_integer(addra);
			douta <= mem(addr_in);
		end if;
	end process;

end RTL;



