library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;

entity prom is

	port (
		clka : in std_logic;
		addra : in std_logic_vector(10 downto 0);
		douta : out std_logic_vector(31 downto 0));

end prom;

architecture RTL of prom is
	subtype word_t is std_logic_vector(31 downto 0);
	type mem_t is array (0 to 2047) of word_t;
	signal addr_in	: integer range 0 to 2047;

	constant mem : mem_t := (
x"00000018",
x"00000000",
x"3f800000",
x"bf800000",
x"00800000",
x"4b000000",
x"4b000000",
x"080001c5",
x"a0000000",
x"a0000000",
x"a0000000",
x"a0630002",
x"a0000000",
x"a0000000",
x"00622820",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"a0000000",
x"68a2000f",
x"a0000000",
x"a0000000",
x"28a2000c",
x"a0000000",
x"a0000000",
x"ac440000",
x"a0000000",
x"a0000000",
x"20420004",
x"a0000000",
x"a0000000",
x"08000014",
x"a0000000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"a0630002",
x"a0000000",
x"a0000000",
x"00622020",
x"a0000000",
x"a0000000",
x"20430000",
x"a0000000",
x"a0000000",
x"a0000000",
x"6882000f",
x"a0000000",
x"a0000000",
x"2882000c",
x"a0000000",
x"a0000000",
x"e4400000",
x"a0000000",
x"a0000000",
x"20420004",
x"a0000000",
x"a0000000",
x"08000032",
x"a0000000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"20030000",
x"c4640000",
x"a0000000",
x"a0000000",
x"e880003d",
x"a0000000",
x"a0000000",
x"c880003a",
x"a0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"20030010",
x"c4620000",
x"a0000000",
x"a0000000",
x"e802000c",
x"a0000000",
x"a0000000",
x"c8020009",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"44200807",
x"a0000000",
x"a0000000",
x"e820004e",
x"a0000000",
x"a0000000",
x"c820004b",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"20030004",
x"c4630000",
x"a0000000",
x"a0000000",
x"44030000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"20030010",
x"c4620000",
x"a0000000",
x"a0000000",
x"e8020009",
x"a0000000",
x"a0000000",
x"c8020006",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"44000806",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"e801000d",
x"a0000000",
x"a0000000",
x"c801000a",
x"a0000000",
x"a0000000",
x"20030004",
x"c4630000",
x"a0000000",
x"a0000000",
x"44030001",
x"a0000000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"c0000046",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"68030012",
x"a0000000",
x"a0000000",
x"2803000f",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"c00000e7",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"20050010",
x"c4a10000",
x"a0000000",
x"a0000000",
x"20050014",
x"8ca40000",
x"a0000000",
x"a0000000",
x"2005000c",
x"8ca50000",
x"a0000000",
x"a0000000",
x"68a30015",
x"a0000000",
x"a0000000",
x"28a30012",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"44010001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040000",
x"c4820000",
x"a0000000",
x"a0000000",
x"a0000000",
x"00651822",
x"a0000000",
x"a0000000",
x"44411000",
x"a0000000",
x"a0000000",
x"68a3fff9",
x"a0000000",
x"a0000000",
x"28a3fff6",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"44010001",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"20030000",
x"c4610000",
x"a0000000",
x"a0000000",
x"e8200012",
x"a0000000",
x"a0000000",
x"c820000f",
x"a0000000",
x"a0000000",
x"44000007",
x"a0000000",
x"a0000000",
x"c0000144",
x"a0000000",
x"a0000000",
x"00031822",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"c0000046",
x"a0000000",
x"a0000000",
x"20040010",
x"c4820000",
x"a0000000",
x"a0000000",
x"20040014",
x"8c840000",
x"a0000000",
x"a0000000",
x"e8400015",
x"a0000000",
x"a0000000",
x"c8400012",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c230000",
x"a0000000",
x"a0000000",
x"00641822",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"2005000c",
x"8ca50000",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"a0000000",
x"44020001",
x"a0000000",
x"a0000000",
x"00651820",
x"a0000000",
x"a0000000",
x"e840fff9",
x"a0000000",
x"a0000000",
x"c840fff6",
x"a0000000",
x"a0000000",
x"44020000",
x"a0000000",
x"a0000000",
x"e4200000",
x"a0000000",
x"a0000000",
x"8c250000",
x"a0000000",
x"a0000000",
x"00a42822",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"0800012d",
x"a0000000",
x"a0000000",
x"a0000000",
x"20030000",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"a0630008",
x"a0000000",
x"a0000000",
x"04002000",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"c0000190",
x"a0000000",
x"a0000000",
x"ac230000",
x"a0000000",
x"a0000000",
x"c4200000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"203f0000",
x"a0000000",
x"a0000000",
x"40210020",
x"a0000000",
x"a0000000",
x"201c0001",
x"a0000000",
x"a0000000",
x"201dffff",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20004",
x"a0000000",
x"a0000000",
x"40210004",
x"a0000000",
x"a0000000",
x"c000000a",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20008",
x"a0000000",
x"a0000000",
x"c000000a",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e2000c",
x"a0000000",
x"a0000000",
x"c000000a",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20010",
x"a0000000",
x"a0000000",
x"c000000a",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040001",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20014",
x"a0000000",
x"a0000000",
x"c000000a",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20030001",
x"a0000000",
x"a0000000",
x"20040000",
x"a0000000",
x"a0000000",
x"afe2001c",
x"a0000000",
x"a0000000",
x"43e20018",
x"a0000000",
x"a0000000",
x"c000000a",
x"a0000000",
x"a0000000",
x"8fe2001c",
x"a0000000",
x"a0000000",
x"20040006",
x"a0000000",
x"a0000000",
x"c00004fc",
x"a0000000",
x"a0000000",
x"20680000",
x"a0000000",
x"a0000000",
x"c0000284",
x"a0000000",
x"a0000000",
x"20210004",
x"a0000000",
x"a0000000",
x"0000003f",
x"a0000000",
x"a0000000",
x"a0000000",
x"00a61820",
x"a0000000",
x"a0000000",
x"a8640001",
x"a0000000",
x"a0000000",
x"00874818",
x"a0000000",
x"a0000000",
x"00c51822",
x"a0000000",
x"a0000000",
x"6b830009",
x"a0000000",
x"a0000000",
x"20a30000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"69280013",
x"a0000000",
x"a0000000",
x"49280009",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"20860000",
x"a0000000",
x"a0000000",
x"08000253",
x"a0000000",
x"a0000000",
x"a0000000",
x"20850000",
x"a0000000",
x"a0000000",
x"08000253",
x"a0000000",
x"a0000000",
x"a0000000",
x"6900026a",
x"a0000000",
x"a0000000",
x"3ce005f5",
x"a0000000",
x"a0000000",
x"1ce0e100",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"20060003",
x"a0000000",
x"a0000000",
x"ac280000",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"3c8005f5",
x"a0000000",
x"a0000000",
x"1c80e100",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280000",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"68030009",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"080002c5",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"3ce00098",
x"a0000000",
x"a0000000",
x"1ce09680",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280004",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"3c800098",
x"a0000000",
x"a0000000",
x"1c809680",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280004",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49400009",
x"a0000000",
x"a0000000",
x"200b0000",
x"a0000000",
x"a0000000",
x"08000306",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"08000317",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"3ce0000f",
x"a0000000",
x"a0000000",
x"1ce04240",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280008",
x"a0000000",
x"a0000000",
x"40210010",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"20210010",
x"a0000000",
x"a0000000",
x"3c80000f",
x"a0000000",
x"a0000000",
x"1c804240",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280008",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49600009",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"08000358",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"08000369",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"3ce00001",
x"a0000000",
x"a0000000",
x"1ce086a0",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac28000c",
x"a0000000",
x"a0000000",
x"40210014",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"20210014",
x"a0000000",
x"a0000000",
x"3c800001",
x"a0000000",
x"a0000000",
x"1c8086a0",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c28000c",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49400009",
x"a0000000",
x"a0000000",
x"200b0000",
x"a0000000",
x"a0000000",
x"080003aa",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"080003bb",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"20072710",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280010",
x"a0000000",
x"a0000000",
x"40210018",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"20210018",
x"a0000000",
x"a0000000",
x"20042710",
x"a0000000",
x"a0000000",
x"00642018",
x"a0000000",
x"a0000000",
x"8c280010",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49600009",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"080003f6",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"08000407",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"200703e8",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280014",
x"a0000000",
x"a0000000",
x"4021001c",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"2021001c",
x"a0000000",
x"a0000000",
x"606403e8",
x"a0000000",
x"a0000000",
x"8c280014",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49400009",
x"a0000000",
x"a0000000",
x"200b0000",
x"a0000000",
x"a0000000",
x"0800043f",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"08000450",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200b0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"20070064",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac280018",
x"a0000000",
x"a0000000",
x"40210020",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"20210020",
x"a0000000",
x"a0000000",
x"60640064",
x"a0000000",
x"a0000000",
x"8c280018",
x"a0000000",
x"a0000000",
x"01044022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49600009",
x"a0000000",
x"a0000000",
x"200a0000",
x"a0000000",
x"a0000000",
x"08000488",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"08000499",
x"a0000000",
x"a0000000",
x"a0000000",
x"20040030",
x"a0000000",
x"a0000000",
x"00831820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"200a0001",
x"a0000000",
x"a0000000",
x"a0000000",
x"2007000a",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"2006000a",
x"a0000000",
x"a0000000",
x"ac28001c",
x"a0000000",
x"a0000000",
x"40210024",
x"a0000000",
x"a0000000",
x"c0000253",
x"a0000000",
x"a0000000",
x"20210024",
x"a0000000",
x"a0000000",
x"6064000a",
x"a0000000",
x"a0000000",
x"8c28001c",
x"a0000000",
x"a0000000",
x"01042022",
x"a0000000",
x"a0000000",
x"6803001d",
x"a0000000",
x"a0000000",
x"49400009",
x"a0000000",
x"a0000000",
x"20050000",
x"a0000000",
x"a0000000",
x"080004d1",
x"a0000000",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20050001",
x"a0000000",
x"a0000000",
x"a0000000",
x"080004e2",
x"a0000000",
x"a0000000",
x"a0000000",
x"20050030",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"20050001",
x"a0000000",
x"a0000000",
x"a0000000",
x"20030030",
x"a0000000",
x"a0000000",
x"00641820",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"2003002d",
x"a0000000",
x"a0000000",
x"04600001",
x"a0000000",
x"a0000000",
x"00084022",
x"a0000000",
x"a0000000",
x"08000284",
x"a0000000",
x"a0000000",
x"a0000000",
x"6b840009",
x"a0000000",
x"a0000000",
x"20830000",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"a0000000",
x"40830001",
x"a0000000",
x"a0000000",
x"ac240000",
x"a0000000",
x"a0000000",
x"20640000",
x"a0000000",
x"a0000000",
x"40210008",
x"a0000000",
x"a0000000",
x"c00004fc",
x"a0000000",
x"a0000000",
x"20210008",
x"a0000000",
x"a0000000",
x"20650000",
x"a0000000",
x"a0000000",
x"8c240000",
x"a0000000",
x"a0000000",
x"40840002",
x"a0000000",
x"a0000000",
x"ac250004",
x"a0000000",
x"a0000000",
x"4021000c",
x"a0000000",
x"a0000000",
x"c00004fc",
x"a0000000",
x"a0000000",
x"2021000c",
x"a0000000",
x"a0000000",
x"8c250004",
x"a0000000",
x"a0000000",
x"00a31820",
x"a0000000",
x"a0000000",
x"e0000000",
x"a0000000",
x"a0000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000"
	 );


begin
	prom_sim: process(clka)
	begin
		if rising_edge(clka) then
			addr_in <= conv_integer(addra);
			douta <= mem(addr_in);
		end if;
	end process;

end RTL;



